`timescale 1ns / 100ps

module sdram_ref_tb;

    logic clk, rst;

    localparam int DATA_WIDTH    = 32;

    localparam real FREQ_MHZ    = 50;
    localparam int ADDR_WIDTH    = 32;
    localparam int SDADDR_WIDTH  = 24;
    localparam int COL_WIDTH     = 9;
    localparam int CAS_LATENCY   = 2;

    parameter DEBUG_SDRAM         = 1;

    localparam real tRC_NS        = 60.0;   // min time in ns between row activations (same bank)
    localparam real tRAS_NS       = 42.0;   // min time in ns from row activation to precharge (same bank)
    localparam real tRCD_NS       = 15.0;   // min time in ns from row activation to read/write
    localparam real tRP_NS        = 15.0;   // min time in ns from precharge to refresh/activation (same bank)
    localparam real tXSR_NS       = 72.0;   // min time in ns from self-refresh exit to activation
    localparam real tREF_NS       = 64e6;   // max time in ns to perform all 8k refresh cycles
    localparam int DELAY_RRD     = 2;       // min clocks between row activations (different bank)
    localparam int DELAY_WR      = 2;       // min clocks write recovery time
    localparam int DELAY_RSC     = 2;       // min clocks for mode register reset

    localparam real CLK_PERIOD=1000/FREQ_MHZ;
    localparam real HALF_CLK_PERIOD=CLK_PERIOD/2;
    localparam real QTR_CLK_PERIOD=CLK_PERIOD/4;
    localparam real OFFSET_CLK_PERIOD=CLK_PERIOD*2/3;
    localparam real IO_LATENCY_NS=CLK_PERIOD/2;
    
    initial
     begin
        $dumpfile("sdram.vcd");
        $dumpvars(0,sdram_core_tb);
        $dumpon;
        #3000000;
        $finish;
     end
    
    initial begin
        clk = 0;
        rst = 1;
        repeat(10) @(posedge clk);
        rst = 0;
    end
    
    always begin
        #HALF_CLK_PERIOD;
        clk = ~clk;
    end
    // clock ram with 90deg lag
    wire #OFFSET_CLK_PERIOD sdram_clk = clk; 

    sdram_ctrl_if #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH)) ctrl_if();
    sdram_dev_if #(.ADDR_WIDTH(SDADDR_WIDTH), .COL_WIDTH(COL_WIDTH)) dev_if();
    
    logic [ADDR_WIDTH-1:0] addr;
    logic [DATA_WIDTH-1:0] read_data, write_data;
    int n;
    always begin
        while(rst) @(posedge clk);
    
        n = 5;
        addr = n<<2;
        write_data = n;

        ctrl_if.addr = addr;
        ctrl_if.write_data = write_data;
        ctrl_if.wr = '1;
        while(~ctrl_if.rdy) @(posedge clk);
        @(posedge clk);
        ctrl_if.wr = '0;
        ctrl_if.write_data = 0;
        while(~ctrl_if.wvalid) @(posedge clk);
        @(posedge clk);
        @(posedge clk);

        ctrl_if.addr = addr;
        ctrl_if.rd = 1;
        while(~ctrl_if.rdy) @(posedge clk);
        @(posedge clk);
        ctrl_if.rd = 0;
        while(~ctrl_if.rvalid) @(posedge clk);
        @(posedge clk);
        @(posedge clk);
        $finish;

        // repeat(1) begin
        //     for (int n = 0; n < 16; n++) begin
        //         addr = n << 10;
        //         write_data = ((n^ 32'hffffffff) << 16) + n;

        //         // write(ctrl_if, clk, addr, write_data);
        //         ctrl_if.addr = addr;
        //         ctrl_if.write_data = write_data;
        //         ctrl_if.wr = '1;
        //         while(~ctrl_if.rdy) @(posedge clk);
        //         @(posedge clk);
        //         ctrl_if.wr = '0;
        //         ctrl_if.write_data = 0;
        //         while(~ctrl_if.wvalid) @(posedge clk);
        //         @(posedge clk);
        //         @(posedge clk);
        //         $display("at time %t Wrote 0x%0x to 0x%0x", $time, write_data, addr);
        //     end            
        //     for (int n = 0; n < 16; n++) begin
        //         addr = n << 10;
        //         write_data = ((n^ 32'hffffffff) << 16) + n;

        //         ctrl_if.addr = addr;
        //         ctrl_if.rd = 1;
        //         while(~ctrl_if.rdy) @(posedge clk);
        //         @(posedge clk);
        //         ctrl_if.rd = 0;
        //         while(~ctrl_if.rvalid) @(posedge clk);
        //         read_data = ctrl_if.read_data;
        //         if(read_data == write_data) $display("at time  %t: Read correct value 0x%0x from 0x%0x", $time, read_data, addr);
        //         else begin
        //             $display("at time %t ERROR: Read incorrect value 0x%0x from 0x%0x, expected 0x%0x", $time, read_data, addr, write_data);
        //             @(posedge clk);
        //             @(posedge clk);
        //             @(posedge clk);
        //             @(posedge clk);
        //             @(posedge clk);
        //             $finish;
        //         end
        //     end            

        // end
        
        // $finish;
    end

    sdram_core_pc
    u_sdram_controller(
        .clk      (clk      ),
        .rst      (rst      ),
        .ctrl_if  (ctrl_if.man),
        .dev_if   (dev_if.sub)
    );

    // spoof ref design to check consistency
    sdram_ctrl_if #(.ADDR_WIDTH(ADDR_WIDTH), .DATA_WIDTH(DATA_WIDTH)) ctrl_if2();
    sdram_dev_if #(.ADDR_WIDTH(SDADDR_WIDTH), .COL_WIDTH(COL_WIDTH)) dev_if2();

    assign ctrl_if2.wr = ctrl_if.wr;
    assign ctrl_if2.rd = ctrl_if.rd;
    assign ctrl_if2.addr = ctrl_if.addr;
    assign ctrl_if2.write_data = ctrl_if.write_data;
    assign dev_if2.read_data = dev_if.read_data;


    wire cmd_diff = dev_if.cmd != dev_if2.cmd;

    sdram_core_ref
    u_sdram_controller_ref(
        .clk      (clk      ),
        .rst      (rst      ),
        .ctrl_if  (ctrl_if2.man),
        .dev_if   (dev_if2.sub)
    );

    

    MT48LC8M16A2 #(
    .IO_LATENCY_NS(IO_LATENCY_NS),
    .Debug(DEBUG_SDRAM),
    .tMRD   (DELAY_RSC*CLK_PERIOD),
    .tRAS   (tRAS_NS),
    .tRC    (tRC_NS),
    .tRCD   (tRCD_NS),
    .tRP    (tRP_NS),
    .tRRD   (DELAY_RRD*CLK_PERIOD)
    )
    u_sdram_model(sdram_clk, dev_if.man);


    // task write(
    //     virtual sdram_ctrl_if ctrl_if,
    //     ref logic  clk,
    //     input logic  [ ADDR_WIDTH-1:0]  a,
    //     input logic  [ DATA_WIDTH-1:0]  data
    //     );

    //     ctrl_if.addr = a;
    //     ctrl_if.write_data = data;
    //     ctrl_if.wr = '1;
    //     while(~ctrl_if.rdy) @(posedge clk);
    //     @(posedge clk);
    //     ctrl_if.wr = '0;
    //     ctrl_if.write_data = 0;
    //     while(~ctrl_if.wvalid) @(posedge clk);
    // endtask

    // task read(
    //     virtual sdram_ctrl_if ctrl_if,
    //     ref logic  clk,
    //     input logic  [ ADDR_WIDTH-1:0]  a,
    //     output logic  [ DATA_WIDTH-1:0]  data
    //     );

    //     ctrl_if.addr = a;
    //     ctrl_if.rd = 1;
    //     while(~ctrl_if.rdy) @(posedge clk);
    //     @(posedge clk);
    //     ctrl_if.rd = 0;
    //     while(~ctrl_if.rvalid) @(posedge clk);
    //     data = ctrl_if.read_data;
    // endtask

endmodule
